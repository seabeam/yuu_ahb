/////////////////////////////////////////////////////////////////////////////////////
// Copyright 2019 seabeam@yahoo.com - Licensed under the Apache License, Version 2.0
// For more information, see LICENCE in the main folder
/////////////////////////////////////////////////////////////////////////////////////
`ifndef YUU_AHB_SLAVE_MEMORY_SV
`define YUU_AHB_SLAVE_MEMORY_SV

typedef yuu_common_memory yuu_ahb_slave_memory;

`endif