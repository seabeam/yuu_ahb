/////////////////////////////////////////////////////////////////////////////////////
// Copyright 2019 seabeam@yahoo.com - Licensed under the Apache License, Version 2.0
// For more information, see LICENCE in the main folder
/////////////////////////////////////////////////////////////////////////////////////
`ifndef YUU_AHB_COMMON_PKG_SVH
`define YUU_AHB_COMMON_PKG_SVH
  
  `include "yuu_ahb_type.sv"
  `include "yuu_ahb_error.sv"
  `include "yuu_ahb_agent_config.sv"
  `include "yuu_ahb_item.sv"

`endif
