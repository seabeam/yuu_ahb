/////////////////////////////////////////////////////////////////////////////////////
// Copyright 2019 seabeam@yahoo.com - Licensed under the Apache License, Version 2.0
// For more information, see LICENCE in the main folder
/////////////////////////////////////////////////////////////////////////////////////
`ifndef YUU_AHB_ENV_PKG_SVH
`define YUU_AHB_ENV_PKG_SVH

  `include "yuu_ahb_env_config.sv"
  `include "yuu_ahb_env.sv"

`endif
