///////////////////////////////////////////////////////////////////////////////////
// Copyright 2019 seabeam@yahoo.com - Licensed under the Apache License, Version 2.0
// For more information, see LICENCE in the main folder
/////////////////////////////////////////////////////////////////////////////////////
`ifndef YUU_AHB_SLAVE_DRIVER_SV
`define YUU_AHB_SLAVE_DRIVER_SV

class yuu_ahb_slave_driver extends uvm_driver #(yuu_ahb_slave_item);
  virtual yuu_ahb_slave_interface  vif;
  uvm_analysis_port #(yuu_ahb_slave_item) out_driver_ap;

  yuu_ahb_slave_config  cfg;
  uvm_event_pool events;

  protected yuu_ahb_slave_memory m_mem;
  
  `uvm_component_utils_begin(yuu_ahb_slave_driver)
  `uvm_component_utils_end

  extern                   function      new(string name, uvm_component parent);
  extern           virtual function void build_phase(uvm_phase phase);
  extern           virtual task          reset_phase(uvm_phase phase);
  extern           virtual task          main_phase(uvm_phase phase);

  extern protected virtual function void init_mem();
  extern protected virtual task          reset_signal();
  extern protected virtual task          get_and_drive();
  extern protected virtual task          drive_bus();
  extern protected virtual task          wait_reset(uvm_phase phase);
endclass

function yuu_ahb_slave_driver::new(string name, uvm_component parent);
  super.new(name, parent);
endfunction

function void yuu_ahb_slave_driver::build_phase(uvm_phase phase);
  out_driver_ap = new("out_driver_ap", this);
  init_mem();
endfunction

task yuu_ahb_slave_driver::reset_phase(uvm_phase phase);
  reset_signal();
endtask

task yuu_ahb_slave_driver::main_phase(uvm_phase phase);
  wait(vif.hreset_n === 1'b1);
  @(vif.cb);
  fork
    get_and_drive();
    wait_reset(phase);
  join
endtask


task yuu_ahb_slave_driver::reset_signal();
  vif.cb.hresp    <= OKAY;
  vif.cb.hready_o <= 1'b1;
  vif.cb.hrdata   <= 'h0;
endtask

function void yuu_ahb_slave_driver::init_mem();
  if (!uvm_config_db #(yuu_ahb_slave_memory)::get(null, get_full_name(), "mem", m_mem))
    m_mem = yuu_ahb_slave_memory::type_id::create("m_mem");
endfunction

task yuu_ahb_slave_driver::get_and_drive();
  forever begin
    drive_bus();
  end
endtask

task yuu_ahb_slave_driver::drive_bus();
  yuu_ahb_addr_t      addr;
  yuu_ahb_direction_e direction;
  yuu_ahb_size_e      size;
  yuu_ahb_data_t      wdata;
  yuu_ahb_data_t      rdata;

  while((vif.cb.htrans !== NONSEQ && vif.cb.htrans !== SEQ) || vif.cb.hsel !== 1'b1 || vif.cb.hready_i !== 1'b1) begin
    @(vif.cb);
  end
  addr = vif.cb.haddr;
  direction = yuu_ahb_direction_e'(vif.cb.hwrite);
  size = yuu_ahb_size_e'(vif.cb.hsize);
  seq_item_port.get_next_item(req); 
  fork
    wait((vif.cb.htrans === NONSEQ || vif.cb.htrans === SEQ) && vif.cb.hsel === 1'b1 && vif.cb.hready_i === 1'b1);
    begin
      vif.cb.hready_o <= 1'b0;
      vif.cb.hresp <= OKAY;
      repeat(req.wait_delay) @(vif.cb);
      if (req.response[0] == ERROR) begin
        vif.cb.hresp <= req.response[0];
        @(vif.cb);
      end
      vif.cb.hready_o <= 1'b1;
    end
  join
  if (direction == WRITE) begin
    yuu_ahb_addr_t low_boundary = addr[7:0] % (`YUU_AHB_ADDR_WIDTH/8);
    yuu_ahb_addr_t high_boundary = low_boundary+(1<<int'(size));
    yuu_ahb_addr_t mem_addr = addr/(`YUU_AHB_ADDR_WIDTH/8);
    int strobe = 0;
    
    for (yuu_ahb_addr_t i=low_boundary; i<high_boundary; i++)
      strobe[i] = 1'b1;

    @(vif.cb);
    wdata = vif.cb.hwdata; 
    vif.cb.hresp <= OKAY;
    if (req.response[0] != ERROR)
      m_mem.write(mem_addr, wdata, strobe);
    seq_item_port.item_done();
  end
  else begin
    yuu_ahb_addr_t mem_addr = addr/(`YUU_AHB_ADDR_WIDTH/8);
    m_mem.read(mem_addr, rdata);
    if (req.response[0] != ERROR)
      if (cfg.use_random_data)
        vif.cb.hrdata <= $urandom();
      else
        vif.cb.hrdata <= rdata;
    else
      vif.cb.hrdata <= 'h0;
    seq_item_port.item_done();
    @(vif.cb);
    vif.cb.hresp <= OKAY;
  end
endtask

task yuu_ahb_slave_driver::wait_reset(uvm_phase phase);
  @(negedge vif.hreset_n);
  phase.jump(uvm_reset_phase::get());
endtask

`endif
