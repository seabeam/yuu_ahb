/////////////////////////////////////////////////////////////////////////////////////
// Copyright 2019 seabeam@yahoo.com - Licensed under the Apache License, Version 2.0
// For more information, see LICENCE in the main folder
/////////////////////////////////////////////////////////////////////////////////////
`ifndef YUU_AHB_MASTER_PKG_SVH
`define YUU_AHB_MASTER_PKG_SVH

  `include "yuu_ahb_master_config.sv"
  `include "yuu_ahb_master_item.sv"
  `include "yuu_ahb_master_sequence_lib.sv"
  `include "yuu_ahb_master_callbacks.sv"
  `include "yuu_ahb_master_driver.sv"
  `include "yuu_ahb_master_monitor.sv"
  `include "yuu_ahb_master_analyzer.sv"
  `include "yuu_ahb_master_collector.sv"
  `include "yuu_ahb_master_adapter.sv"
  `include "yuu_ahb_master_agent.sv"

`endif
